--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   23:53:32 04/24/2016
-- Design Name:   
-- Module Name:   C:/Users/Angela/Desktop/oscar/arquitectura/procesadorIII/SEU_tb.vhd
-- Project Name:  procesadorIII
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: SEU
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY SEU_tb IS
END SEU_tb;
 
ARCHITECTURE behavior OF SEU_tb IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT SEU
    PORT(
         EntradaSEU : IN  std_logic_vector(12 downto 0);
         SalidaSEU : OUT  std_logic_vector(31 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal EntradaSEU : std_logic_vector(12 downto 0) := (others => '0');

 	--Outputs
   signal SalidaSEU : std_logic_vector(31 downto 0);
   -- No clocks detected in port list. Replace <clock> below with 
   -- appropriate port name 
 
  
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: SEU PORT MAP (
          EntradaSEU => EntradaSEU,
          SalidaSEU => SalidaSEU
        );

   --
 

   -- Stimulus process
   stim_proc: process
   begin		
--      EntradaSEU <= "0000000000110";
--		wait for 100 ns;
--		EntradaSEU <= "1000000000110"; 
		
  --    wait;
   end process;

END;